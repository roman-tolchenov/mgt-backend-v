module mgt

fn test_event() {
    assert true
}
