module main
import mgt

fn main() {
    println('Hello World! ${mgt.a}')
}
